mi_pll_divisor_inst : mi_pll_divisor PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
