pll_dividerx2_inst : pll_dividerx2 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
